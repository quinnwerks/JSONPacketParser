`timescale 1 ns/ 1ps

// Struct for flit data
 typedef struct packed {
    int data;
    int keep;
    int last;
} flit;

// Struct for packet data (max 23 flits)
typedef struct packed {
    flit [22:0] flit_list;
    int num_flits;
} packet;

// DPI
import "DPI-C" function packet parseJSON(input string jsonFilePath, input int ver);

// Top
module testbench();

    reg clk;
    reg resetn;
    
    reg [7:0] keep;
    reg last;
    reg [63:0] data;
    reg valid;
    
    wire ready;
 
    reg ready_reg;
    reg ready_out;
    
    wire [2:0] state;
    wire state_valid;
    
    always #5 clk = ~clk;
    
    always@(posedge clk)
    begin
        ready_reg <= ready;
    end
    
    initial begin
        ready_out = 1;
        clk = 0;
        #5 resetn = 1;
    end

    initial begin
        string jsonFilePath = "../jsonTests/jsonPacketTest_extensive.json";
        int ver = 1'd0;
        packet [63:0] packetList = parseJSON(jsonFilePath, ver);
    end

    initial begin
        #50

        gen_transaction(64'd0, 64'hc4c0c02ca553e16fa, 8'hff, 1'b0);
        gen_transaction(64'd1, 64'h0000007447c0887a, 8'hff, 1'b0);
        gen_transaction(64'd2, 64'h0100000100030000, 8'hff, 1'b0);
        gen_transaction(64'd3, 64'h5073930200000000, 8'h0f, 1'b1);
    end
    
wire [63:0] data_out;
wire [7:0] keep_out;
wire last_out;
wire valid_out;

wire [47:0] observedAddress_out;
wire observedAddress_out_valid;

/*
design_1 design_1_i
   (.M_AXIS_tdata(data_out),
    .M_AXIS_tdest(),
    .M_AXIS_tkeep(keep_out),
    .M_AXIS_tlast(last_out),
    .M_AXIS_tready(ready_out),
    .M_AXIS_tvalid(valid_out),
    .S_AXIS_tdata(data),
    .S_AXIS_tkeep(keep),
    .S_AXIS_tlast(last),
    .S_AXIS_tready(ready),
    .S_AXIS_tvalid(valid),
    .aclk_0(clk),
    .aresetn_0(resetn),
    .mac_addr_V_0(48'hfa163e55ca02),
    .observedAddress_out_V_0(observedAddress_out),
    .observedAddress_out_V_ap_vld_0(observedAddress_out_valid),
    .state_out_V_0(state),
    .state_out_V_ap_vld_0(state_valid)
    
    );
   
*/

   pr pr_i
       (.ARESETN(resetn),
        .CLK(clk),
        .M_AXIS_tdata(data_out),
        .M_AXIS_tkeep(keep_out),
        .M_AXIS_tlast(last_out),
        .M_AXIS_tready(ready_out),
        .M_AXIS_tvalid(valid_out),
        .S_AXIS_tdata(data),
        .S_AXIS_tkeep(keep),
        .S_AXIS_tlast(last),
        .S_AXIS_tready(ready),
        .S_AXIS_tvalid(valid),
        .S_AXI_CONTROL_araddr(M_AXI_CONTROL_araddr),
        //.S_AXI_CONTROL_arprot(M_AXI_CONTROL_arprot),
        //.S_AXI_CONTROL_arqos(M_AXI_CONTROL_arqos),
        .S_AXI_CONTROL_arready(M_AXI_CONTROL_arready),
        .S_AXI_CONTROL_arvalid(M_AXI_CONTROL_arvalid),
        .S_AXI_CONTROL_awaddr(M_AXI_CONTROL_awaddr),
        //.S_AXI_CONTROL_awprot(M_AXI_CONTROL_awprot),
        //.S_AXI_CONTROL_awqos(M_AXI_CONTROL_awqos),
        .S_AXI_CONTROL_awready(M_AXI_CONTROL_awready),
        .S_AXI_CONTROL_awvalid(M_AXI_CONTROL_awvalid),
        .S_AXI_CONTROL_bready(M_AXI_CONTROL_bready),
        .S_AXI_CONTROL_bresp(M_AXI_CONTROL_bresp),
        .S_AXI_CONTROL_bvalid(M_AXI_CONTROL_bvalid),
        .S_AXI_CONTROL_rdata(M_AXI_CONTROL_rdata),
        .S_AXI_CONTROL_rready(M_AXI_CONTROL_rready),
        .S_AXI_CONTROL_rresp(M_AXI_CONTROL_rresp),
        .S_AXI_CONTROL_rvalid(M_AXI_CONTROL_rvalid),
        .S_AXI_CONTROL_wdata(M_AXI_CONTROL_wdata),
        .S_AXI_CONTROL_wready(M_AXI_CONTROL_wready),
        .S_AXI_CONTROL_wstrb(M_AXI_CONTROL_wstrb),
        .S_AXI_CONTROL_wvalid(M_AXI_CONTROL_wvalid),
        .S_AXI_MEM_0_araddr(S_AXI_MEM_0_araddr),
        .S_AXI_MEM_0_arburst(S_AXI_MEM_0_arburst),
        .S_AXI_MEM_0_arcache(S_AXI_MEM_0_arcache),
        //.S_AXI_MEM_0_arid(S_AXI_MEM_0_arid),
        .S_AXI_MEM_0_arlen(S_AXI_MEM_0_arlen),
        .S_AXI_MEM_0_arlock(S_AXI_MEM_0_arlock),
        .S_AXI_MEM_0_arprot(S_AXI_MEM_0_arprot),
        .S_AXI_MEM_0_arqos(S_AXI_MEM_0_arqos),
        .S_AXI_MEM_0_arready(S_AXI_MEM_0_arready),
        .S_AXI_MEM_0_arsize(S_AXI_MEM_0_arsize),
        .S_AXI_MEM_0_arvalid(S_AXI_MEM_0_arvalid),
        .S_AXI_MEM_0_awaddr(S_AXI_MEM_0_awaddr),
        .S_AXI_MEM_0_awburst(S_AXI_MEM_0_awburst),
        .S_AXI_MEM_0_awcache(S_AXI_MEM_0_awcache),
        //.S_AXI_MEM_0_awid(S_AXI_MEM_0_awid),
        .S_AXI_MEM_0_awlen(S_AXI_MEM_0_awlen),
        .S_AXI_MEM_0_awlock(S_AXI_MEM_0_awlock),
        .S_AXI_MEM_0_awprot(S_AXI_MEM_0_awprot),
        .S_AXI_MEM_0_awqos(S_AXI_MEM_0_awqos),
        .S_AXI_MEM_0_awready(S_AXI_MEM_0_awready),
        .S_AXI_MEM_0_awsize(S_AXI_MEM_0_awsize),
        .S_AXI_MEM_0_awvalid(S_AXI_MEM_0_awvalid),
        //.S_AXI_MEM_0_bid(S_AXI_MEM_0_bid),
        .S_AXI_MEM_0_bready(S_AXI_MEM_0_bready),
        .S_AXI_MEM_0_bresp(S_AXI_MEM_0_bresp),
        .S_AXI_MEM_0_bvalid(S_AXI_MEM_0_bvalid),
        .S_AXI_MEM_0_rdata(S_AXI_MEM_0_rdata),
        //.S_AXI_MEM_0_rid(S_AXI_MEM_0_rid),
        .S_AXI_MEM_0_rlast(S_AXI_MEM_0_rlast),
        .S_AXI_MEM_0_rready(S_AXI_MEM_0_rready),
        .S_AXI_MEM_0_rresp(S_AXI_MEM_0_rresp),
        .S_AXI_MEM_0_rvalid(S_AXI_MEM_0_rvalid),
        .S_AXI_MEM_0_wdata(S_AXI_MEM_0_wdata),
        .S_AXI_MEM_0_wlast(S_AXI_MEM_0_wlast),
        .S_AXI_MEM_0_wready(S_AXI_MEM_0_wready),
        .S_AXI_MEM_0_wstrb(S_AXI_MEM_0_wstrb),
        .S_AXI_MEM_0_wvalid(S_AXI_MEM_0_wvalid),
        .S_AXI_MEM_1_araddr(S_AXI_MEM_1_araddr),
        .S_AXI_MEM_1_arburst(S_AXI_MEM_1_arburst),
        .S_AXI_MEM_1_arcache(S_AXI_MEM_1_arcache),
        //.S_AXI_MEM_1_arid(S_AXI_MEM_1_arid),
        .S_AXI_MEM_1_arlen(S_AXI_MEM_1_arlen),
        .S_AXI_MEM_1_arlock(S_AXI_MEM_1_arlock),
        .S_AXI_MEM_1_arprot(S_AXI_MEM_1_arprot),
        .S_AXI_MEM_1_arqos(S_AXI_MEM_1_arqos),
        .S_AXI_MEM_1_arready(S_AXI_MEM_1_arready),
        .S_AXI_MEM_1_arsize(S_AXI_MEM_1_arsize),
        .S_AXI_MEM_1_arvalid(S_AXI_MEM_1_arvalid),
        .S_AXI_MEM_1_awaddr(S_AXI_MEM_1_awaddr),
        .S_AXI_MEM_1_awburst(S_AXI_MEM_1_awburst),
        .S_AXI_MEM_1_awcache(S_AXI_MEM_1_awcache),
        //.S_AXI_MEM_1_awid(S_AXI_MEM_1_awid),
        .S_AXI_MEM_1_awlen(S_AXI_MEM_1_awlen),
        .S_AXI_MEM_1_awlock(S_AXI_MEM_1_awlock),
        .S_AXI_MEM_1_awprot(S_AXI_MEM_1_awprot),
        .S_AXI_MEM_1_awqos(S_AXI_MEM_1_awqos),
        .S_AXI_MEM_1_awready(S_AXI_MEM_1_awready),
        .S_AXI_MEM_1_awsize(S_AXI_MEM_1_awsize),
        .S_AXI_MEM_1_awvalid(S_AXI_MEM_1_awvalid),
        //.S_AXI_MEM_1_bid(S_AXI_MEM_1_bid),
        .S_AXI_MEM_1_bready(S_AXI_MEM_1_bready),
        .S_AXI_MEM_1_bresp(S_AXI_MEM_1_bresp),
        .S_AXI_MEM_1_bvalid(S_AXI_MEM_1_bvalid),
        .S_AXI_MEM_1_rdata(S_AXI_MEM_1_rdata),
        //.S_AXI_MEM_1_rid(S_AXI_MEM_1_rid),
        .S_AXI_MEM_1_rlast(S_AXI_MEM_1_rlast),
        .S_AXI_MEM_1_rready(S_AXI_MEM_1_rready),
        .S_AXI_MEM_1_rresp(S_AXI_MEM_1_rresp),
        .S_AXI_MEM_1_rvalid(S_AXI_MEM_1_rvalid),
        .S_AXI_MEM_1_wdata(S_AXI_MEM_1_wdata),
        .S_AXI_MEM_1_wlast(S_AXI_MEM_1_wlast),
        .S_AXI_MEM_1_wready(S_AXI_MEM_1_wready),
        .S_AXI_MEM_1_wstrb(S_AXI_MEM_1_wstrb),
        .S_AXI_MEM_1_wvalid(S_AXI_MEM_1_wvalid)
    );

// Get transaction task
task gen_transaction(input [63:0] num, input [63:0] data_task, input [7:0] keep_task, input last_task);

  data = data_task;
  keep = keep_task;
  last = last_task;
  wait(ready);
  valid = 1;
  #10
  $display("Transaction %d, Data: %h, keep %h, last %b", num, data_task, keep_task, last_task);
  
endtask

endmodule